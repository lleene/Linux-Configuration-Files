VERSION 5.5 ;
UNITS
    CURRENT MILLIAMPS 10000 ;
    VOLTAGE VOLTS 1000 ;
    FREQUENCY MEGAHERTZ 10 ;
    CAPACITANCE PICOFARADS 10 ;
    DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

LAYER POLY1
    TYPE MASTERSLICE ;
END POLY1
